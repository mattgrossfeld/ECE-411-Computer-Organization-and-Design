library verilog;
use verilog.vl_types.all;
entity cache_L2_4way_control is
    port(
        counter_pick    : out    vl_logic_vector(1 downto 0);
        clk             : in     vl_logic;
        hit_sel         : out    vl_logic_vector(1 downto 0);
        hit0            : in     vl_logic;
        hit1            : in     vl_logic;
        hit2            : in     vl_logic;
        hit3            : in     vl_logic;
        write_data0     : out    vl_logic;
        write_data1     : out    vl_logic;
        write_data2     : out    vl_logic;
        write_data3     : out    vl_logic;
        write_tag0      : out    vl_logic;
        write_tag1      : out    vl_logic;
        write_tag2      : out    vl_logic;
        write_tag3      : out    vl_logic;
        write_dirty0    : out    vl_logic;
        write_dirty1    : out    vl_logic;
        write_dirty2    : out    vl_logic;
        write_dirty3    : out    vl_logic;
        write_valid0    : out    vl_logic;
        write_valid1    : out    vl_logic;
        write_valid2    : out    vl_logic;
        write_valid3    : out    vl_logic;
        write_lru       : out    vl_logic;
        valid0          : in     vl_logic;
        valid1          : in     vl_logic;
        valid2          : in     vl_logic;
        valid3          : in     vl_logic;
        valid0_out      : out    vl_logic;
        valid1_out      : out    vl_logic;
        valid2_out      : out    vl_logic;
        valid3_out      : out    vl_logic;
        dirty0          : in     vl_logic;
        dirty1          : in     vl_logic;
        dirty2          : in     vl_logic;
        dirty3          : in     vl_logic;
        dirty0_out      : out    vl_logic;
        dirty1_out      : out    vl_logic;
        dirty2_out      : out    vl_logic;
        dirty3_out      : out    vl_logic;
        lru             : in     vl_logic_vector(2 downto 0);
        lru_out         : out    vl_logic_vector(2 downto 0);
        addr_mux_sel    : out    vl_logic_vector(2 downto 0);
        datainmux_sel   : out    vl_logic;
        mem_read        : in     vl_logic;
        mem_write       : in     vl_logic;
        mem_resp        : out    vl_logic;
        pmem_resp       : in     vl_logic;
        pmem_read       : out    vl_logic;
        pmem_write      : out    vl_logic
    );
end cache_L2_4way_control;
