library verilog;
use verilog.vl_types.all;
entity ewb_sv_unit is
end ewb_sv_unit;
