library verilog;
use verilog.vl_types.all;
entity ewb_control_sv_unit is
end ewb_control_sv_unit;
