library verilog;
use verilog.vl_types.all;
entity pipe_datapath_sv_unit is
end pipe_datapath_sv_unit;
