library verilog;
use verilog.vl_types.all;
entity fwd_logic_sv_unit is
end fwd_logic_sv_unit;
