library verilog;
use verilog.vl_types.all;
entity cache_L2_4way_sv_unit is
end cache_L2_4way_sv_unit;
