library verilog;
use verilog.vl_types.all;
entity cc_comp_sv_unit is
end cc_comp_sv_unit;
