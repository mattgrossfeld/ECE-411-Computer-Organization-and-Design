library verilog;
use verilog.vl_types.all;
entity data_decoder_sv_unit is
end data_decoder_sv_unit;
