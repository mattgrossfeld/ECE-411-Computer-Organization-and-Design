library verilog;
use verilog.vl_types.all;
entity mem_wb_sv_unit is
end mem_wb_sv_unit;
