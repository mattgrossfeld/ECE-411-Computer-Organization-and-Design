library verilog;
use verilog.vl_types.all;
entity ewb_datapath_sv_unit is
end ewb_datapath_sv_unit;
