import rv32i_types::*;

module mp1
(
    input clk,

    /* Memory signals */
    input mem_resp,
    input [31:0] mem_rdata,
    output mem_read,
    output mem_write,
    output [3:0] mem_byte_enable,
    output [31:0] mem_address,
    output [31:0] mem_wdata
);

rv32i_opcode opcode;
logic [2:0] funct3;
logic [6:0] funct7;
//logic bit30;
logic br_en;
logic load_pc;
logic load_ir;
logic load_regfile;
logic load_mar;
logic load_mdr;
logic [1:0] pcmux_sel;
logic [2:0] regfilemux_sel;
logic [1:0] memdatamux_sel;
logic marmux_sel;
alu_ops aluop;
logic alumux1_sel;
logic [2:0] alumux2_sel;
logic addrmux_sel;
branch_funct3_t cmpop;
logic cmpmux_sel;
logic load_data_out;
logic jalr;


/* Instantiate MP 0 top level blocks here */

control control
(
    .clk(clk),
	/* Datapath controls */
	.opcode(opcode),
	.funct3(funct3),
	.funct7(funct7),
//	.bit30(bit30),
	.br_en(br_en),
	.load_pc(load_pc),
	.load_ir(load_ir),
	.load_regfile(load_regfile),
	.load_mar(load_mar),
	.load_mdr(load_mdr),
	.load_data_out(load_data_out),
	.pcmux_sel(pcmux_sel),
	.regfilemux_sel(regfilemux_sel),
	.marmux_sel(marmux_sel),
	.cmpmux_sel(cmpmux_sel),
	.alumux1_sel(alumux1_sel),
	.memdatamux_sel(memdatamux_sel),
	.alumux2_sel(alumux2_sel),
	.aluop(aluop),
	.cmpop(cmpop),
	.mem_resp(mem_resp),
	.mem_read(mem_read),
	.mem_write(mem_write),
	.mem_byte_enable(mem_byte_enable)
);

datapath datapath
(
	.clk(clk),
	.pcmux_sel(pcmux_sel),
	.load_pc(load_pc),
	.cmpmux_sel(cmpmux_sel),
	.load_ir(load_ir),
	.load_regfile(load_regfile),
	.load_mar(load_mar),
	.load_mdr(load_mdr),
	.load_data_out(load_data_out),
	.alumux1_sel(alumux1_sel),
	.alumux2_sel(alumux2_sel),
	.regfilemux_sel(regfilemux_sel),
	.marmux_sel(marmux_sel),
	.aluop(aluop),
	.mem_rdata(mem_rdata),
	.cmpop(cmpop),
	.mem_address(mem_address),
	.mem_wdata(mem_wdata),
	.opcode(opcode),
	.funct3(funct3),
	.memdatamux_sel(memdatamux_sel),
	.funct7(funct7),
//	.bit30(bit30),
	.br_en(br_en)
);

endmodule : mp1
