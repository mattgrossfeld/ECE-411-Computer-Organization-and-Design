library verilog;
use verilog.vl_types.all;
entity stall_load_control_sv_unit is
end stall_load_control_sv_unit;
